class bridge_rbase_seq extends uvm_sequence#(read_xtn);
    `uvm_object_utils(bridge_rbase_seq);
extern function new(string name ="bridge_rbase_seq");
 //extern task body();

endclass
	function bridge_rbase_seq::new(string name ="bridge_rbase_seq");
		super.new(name);
	endfunction
////////////////////////////////////////////////////


